library IEEE;
    use IEEE.std_logic_1164.all;
    use IEEE.numeric_std.all;

entity simple_cpu_tb is
end simple_cpu_tb;

architecture beh of simple_cpu_tb is
    constant clk_period : time := 100 ns;
    constant T_RESET : time := 250 ns;
    constant N          : positive := 8;
    constant M          : positive := 4;

    component simple_cpu is
        generic(
            N : natural := 8; -- number of bits of the registers
            M : natural := 4 -- number of bits of the memory addresses
        );
        port(
            clk : in std_logic;
            rst : in std_logic;
            instr : in std_logic_vector(N-1 downto 0);
            pc : out std_logic_vector(M-1 downto 0);
            input : in std_logic_vector(N-1 downto 0);
            output : out std_logic_vector(N-1 downto 0)
        );
    end component;
    
    signal clk : std_logic := '0';
    signal rst_ext   : std_logic := '0';
    signal instr_ext : std_logic_vector(N-1 downto 0) := (others => '0');
    signal pc_ext : std_logic_vector(M - 1 downto 0);
    signal input_ext : std_logic_vector(N - 1 downto 0) := (others => '0');
    signal output_ext : std_logic_vector(N - 1 downto 0);
    signal testing : boolean := true;
begin

    clk <= not clk after clk_period/2 when testing else '0';
    rst_ext <= '1' after T_RESET;
    
    DUT: simple_cpu
        generic map(
            N => N,
            M => M
        )
        port map (
            clk => clk,
            rst => rst_ext,
            instr => instr_ext,
            pc => pc_ext,
            input => input_ext,
            output => output_ext 
        );

    STIMULI : process(clk, rst_ext)
        variable t : integer := 0;
    begin
        if rst_ext = '0' then
            input_ext <= (others => '0');
            --output_ext <= (others => '0'); -- poi si vedrà 
            instr_ext <= (others => '0');
            --pc_ext <= (others => '0');
            t := 0;
        elsif rising_edge(clk) then
            case t is
                when 0 =>
                when 1 => input_ext <= "00000100";
                when 2 =>
                when 3 =>
                when 4 =>
                when 5 =>
                when 6 =>
                when 7 =>
                when 8 =>
                
                when 25 => testing <= false;
                when others =>
            end case;
            t := t+1;
        end if;
    end process;

end architecture;